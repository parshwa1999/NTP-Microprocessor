`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:04:09 09/01/2017 
// Design Name: 
// Module Name:    Write_Back_Block 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Write_Back_Block(
    output reg [7:0] ans_wb,
    input [7:0] ans_dm,
    input clk,
    input reset
    );
	 
///////////////////////////////////////////////////////////////////////////////////Declarations/////////////////////////////////////////////////////////////////////////////////////////
	 wire[7:0] ans_wb_temp;
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	 
//////////////////////////////////////////////////////////////////////////////////Combinational Block//////////////////////////////////////////////////////////////////////////////////////////// 
	 assign ans_wb_temp = (reset == 1'b0) ? 8'b0000_0000 : ans_dm; // Value to be scanned at next clock edge
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	 
//////////////////////////////////////////////////////////////////////////////////Sequential Block//////////////////////////////////////////////////////////////////////////////////////
	always@(posedge clk)
	begin
		ans_wb <= ans_wb_temp;	// Scanning the value at positive clock edge
	end
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
endmodule
