`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:01:15 08/18/2017 
// Design Name: 
// Module Name:    Data_Memory_Block 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Data_Memory_Block(
	 output [7:0] ans_dm,
    input [7:0] ans_ex,
    input [7:0] DM_data,
    input mem_rw_ex,
    input mem_en_ex,
    input mem_mux_sel_dm,
    input reset,
    input clk
    );
////////////////////////////////////////////////Declartions//////////////////////////////////////////////////////////////////////
	wire [7:0] DM_out, Ex_out_tmp;
	reg [7:0] Ex_out;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////Data Memory Block////////////////////////////////////////////////////////////////
	Data_Memory DM1 (
  .clka(clk), // input clk
  .ena(mem_en_ex), // input mem_en_ex
  .wea(mem_rw_ex), // input [0 : 0] mem_rw_ex
  .addra(ans_ex), // input [7 : 0] ans_ex
  .dina(DM_data), // input [7 : 0] DM_data
  .douta(DM_out) // output [7 : 0] DM_out
);
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	

////////////////////////////////////////////////Combinational Block//////////////////////////////////////////////////////////////
	assign ans_dm = (mem_mux_sel_dm) ? DM_out : Ex_out;	// Mux used as select line
	assign Ex_out_tmp = reset ?  ans_ex : 8'b0000_0000;
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////Sequential Block//////////////////////////////////////////////////////////////////
	always @(posedge clk)
	begin
		Ex_out <= Ex_out_tmp;
	end
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
endmodule