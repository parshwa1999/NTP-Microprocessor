`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:31:57 08/18/2017 
// Design Name: 
// Module Name:    Register_Bank_Block 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Register_Bank_Block(
	output [7:0] A,
    output [7:0] B,
    input [23:0] ins,
    input [7:0] ans_ex,
    input [7:0] ans_dm,
    input [7:0] ans_wb,
    input [7:0] imm,
    input [4:0] RW_dm,
    input [1:0] mux_sel_A,
    input [1:0] mux_sel_B,
    input imm_sel,
    input clk
    );
////////////////////////////////////////////////Declartions//////////////////////////////////////////////////////////////////////	 
	wire [7:0] BI; 
	reg [7:0] reg_bank[0:31];		// Register bank of 8 bits
	reg [7:0] AR, BR;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////Combinational Block//////////////////////////////////////////////////////////////
	assign A = mux_sel_A[0] & mux_sel_A[1] ? ans_wb : mux_sel_A[0] & ~mux_sel_A[1] ? ans_ex : ~mux_sel_A[0] & mux_sel_A[1] ? ans_dm : AR;
	assign BI = mux_sel_B[0] & mux_sel_B[1] ? ans_wb : mux_sel_B[0] & ~mux_sel_B[1] ? ans_ex : ~mux_sel_B[0] & mux_sel_B[1] ? ans_dm : BR;
	assign B = imm_sel ? imm : BI;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
////////////////////////////////////////////////Sequential block/////////////////////////////////////////////////////////////////	
	always@(posedge clk)
	begin
		AR <= reg_bank[ins[13:9]];
		BR <= reg_bank[ins[8:4]];
		reg_bank[RW_dm] <= ans_dm;
	end
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
endmodule
