`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:08:29 08/11/2017 
// Design Name: 
// Module Name:    PCIM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PCIM(
    output [23:0] ins,
    output [7:0] Current_Address,
	 input [7:0] jmp_loc,
    input pc_mux_sel,
    input Stall,
    input Stall_pm,
    input reset,
    input clk
    );

/////////////////////////////////////////////////////////Declarations/////////////////////////////////////////////////////////////////////////////////////////////////////
	wire [7:0] CAJ, CAR, Hold_Address_temp, Next_Address_temp;
	wire [23:0] PM_out, ins_pm;
	wire [23:0] ins_prv_temp;
	
	reg [7:0] Hold_Address, Next_Address;
	reg [23:0] ins_prv;
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////Program Memory//////////////////////////////////////////////////////////////////////////////////////////////////
	Program_Memory pm1(
  .clka(clk), 					// input clk
  .addra(Current_Address), // input [7 : 0] Current_Address
  .douta(PM_out) 				// output [23 : 0] PM_out
	);
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	


//////////////////////////////////////////////////////////////////////////////Combinational block//////////////////////////////////////////////////////////////////////////////////////////////
	assign CAJ = (Stall) ? Hold_Address : Next_Address;
	assign CAR = (pc_mux_sel) ? jmp_loc : CAJ;
	assign Current_Address = (reset) ? CAR : 8'b0000_0000;
	
	assign ins_pm = (Stall_pm) ? ins_prv : PM_out;
	assign ins = (reset) ? ins_pm : 24'b0000_0000_0000_0000_0000_0000;
	
	assign ins_prv_temp = (reset) ? ins : 24'b0000_0000_0000_0000_0000_0000;
	assign Hold_Address_temp = (reset) ? Current_Address : 8'b0000_0000;
	assign Next_Address_temp = (reset) ? Current_Address + 8'b0000_0001 : 8'b0000_0000;
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
//////////////////////////////////////////////////////////////////////////////Sequential block////////////////////////////////////////////////////////////////////////////////////////////////	
	always @ (posedge clk)
	begin
		ins_prv <= ins_prv_temp;
		Hold_Address <= Hold_Address_temp;
		Next_Address <= Next_Address_temp;
	end
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


endmodule
